LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY tb_i2c_esclavo_completo IS
END tb_i2c_esclavo_completo;

ARCHITECTURE behavior OF tb_i2c_esclavo_completo IS

    -- Component declaration of the design under test (DUT)
    COMPONENT i2c_esclavo_completo
        PORT(
            SDA : IN std_logic;
            SCL : IN std_logic;
            reset : IN std_logic;
            SDA_int : OUT std_logic
        );
    END COMPONENT;

    -- Signals to connect to the DUT
    signal SDA     : std_logic := '0';
    signal SCL     : std_logic := '0';
    signal reset   : std_logic := '0';
    signal SDA_int : std_logic;

    -- Clock period definition
    constant clk_period : time := 10 ns;

    -- Vector for SDA sequence (24 bits)
    signal SDA_sequence : std_logic_vector(23 downto 0) := "100100011000100000110000";  

BEGIN

    -- Instantiate the Unit Under Test (UUT)
    uut: i2c_esclavo_completo
        PORT MAP(
            SDA => SDA,
            SCL => SCL,
            reset => reset,
            SDA_int => SDA_int
        );

    -- Clock generation process
    clk_process :process
    begin
        SCL <= '0';
        wait for clk_period / 2;
        SCL <= '1';
        wait for clk_period / 2;
    end process;

    -- Stimulus process
    stim_proc: process
    begin
        -- Reset
        reset <= '1';
        wait for 20 ns;
        reset <= '0';

        -- Wait for the clock to stabilize
        wait for 10 ns;

        -- Inserto SDA
        for i in 0 to 23 loop
            if i = 0 then
                -- Before the first falling edge of SCL, set SDA = 0 (CONDICION DE START)
                SDA <= '0';
                wait until SCL = '1';  -- Wait for the rising edge of SCL
            else
                -- Apply the SDA sequence on the falling edge of SCL
                wait until SCL = '0';  -- Wait for the falling edge of SCL
                SDA <= SDA_sequence(i);
            end if;
        end loop;

        -- Finish simulation after the sequence
        wait for 100 ns;
        assert false report "End of testbench" severity note;
        wait;
    end process;

END behavior;
